module comparator (A,B,F);
input [2:0] A,B;
output F;

assign F=A>B;

    
endmodule